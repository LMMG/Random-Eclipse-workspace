death-signs: true
diamond-ore-notifications: true
death-lightning: true
map-number: 1
kit-map: false
prevent-ally-damage: true
exp-multiplier:
  global: 2.0
  fishing: 2.0
  smelting: 2.0
  looting-per-level: 1.5
  luck-per-level: 1.5
  fortune-per-level: 1.5
roads:
  allow-claims-besides: true
combatlog:
  enabled: true
  despawn-delay-ticks: 600
conquest:
  point-loss-per-death: 20
  victory-points: 300
  allow-negative-points: true
warzone:
  radius: 800
factions:
  disallowed-faction-names:
  - EOTW
  min-name-characters: 3
  max-name-characters: 16
  max-members: 25
  max-allies: 1
subclaims:
  min-name-characters: 3
  max-name-characters: 16
relation-colours:
  wilderness: DARK_GREEN
  warzone: LIGHT_PURPLE
  teammate: GREEN
  ally: GOLD
  enemy: RED
  road: GOLD
deaths-till-raidable:
  maximum: 6
  millis-between-updates: 45000
  increment-between-updates: 0.1
deathban:
  base-duration-minutes: 120
  respawn-screen-seconds-before-kick: 15
enchantment-limits:
  PROTECTION_ENVIRONMENTAL: 3
  PROTECTION_FIRE: 3
  SILK_TOUCH: 1
  DURABILITY: 3
  PROTECTION_EXPLOSIONS: 3
  LOOT_BONUS_BLOCKS: 3
  PROTECTION_PROJECTILE: 3
  OXYGEN: 3
  WATER_WORKER: 1
  THORNS: 0
  DAMAGE_ALL: 3
  ARROW_KNOCKBACK: 1
  KNOCKBACK: 1
  FIRE_ASPECT: 1
  LOOT_BONUS_MOBS: 3
  LUCK: 3
  LURE: 3
end:
  open: true
  exit: world,0.5,75,0.5,0,0
eotw:
  chat-symbol-prefix: ""
  chat-symbol-suffix: ""
  last-map-cappers: []
potion-limits:
  STRENGTH: 0
  INVISIBILITY: 0
  REGEN: 0
  WEAKNESS: 0
  INSTANT_DAMAGE: 0
  SLOWNESS: 1
  POISON: 1
